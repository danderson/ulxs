package ISA

typedef 16 W;

typedef Bit#(W) PC;
typedef Bit#(W) GPR;
typedef Bit#(4) JumpOffset;

endpackage
