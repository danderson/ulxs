package TB;

import Strobe::*;
import StmtFSM::*;

module mkTB ();
   mkStrobeTest();
endmodule

endpackage
